module ShiftLeft2_26to28(input [25:0] IN,output [27:0] S);

	assign S = IN<<2;
	
endmodule