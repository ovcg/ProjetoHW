module ShiftLeft2(input [31:00] IN, output [31:0] S);

	assign S = IN<<2;
	
endmodule